/**
 * @file RegFile.sv
 * @author Jacob Chisholm (https://Jchisholm204.github.io)
 * @brief 
 * @version 0.1
 * @date Created: 2025-05-14
 * @modified Last Modified: 2025-05-14
 *
 * @copyright Copyright (c) 2025
 */

module RegFile(

);

endmodule
