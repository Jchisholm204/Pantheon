/**
 * @file DCSRs.sv
 * @author Jacob Chisholm (https://Jchisholm204.github.io)
 * @brief Debug CSRs
 * @version 0.1
 * @date Created: 2025-08-03
 * @modified Last Modified: 2025-08-03
 *
 * @copyright Copyright (c) 2025
 */

`timescale 1ns/100ps
module DCSRs(
    input logic iClk, nRst
);

endmodule

